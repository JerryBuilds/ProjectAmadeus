`include "Defines.v"

module MusicGenerateFragment (
  input clk, reset,
  
  output done
);