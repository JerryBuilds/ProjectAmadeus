`include "Defines.v"

module MusicFragmentDecomposition (
  input clk, reset,
  
  output done
);