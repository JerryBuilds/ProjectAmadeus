`include "Defines.v"

module MusicMergeFragments (
  input clk, reset,
  
  output done
);